library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;

entity T_Box_2_port is
    port ( CLK : IN  std_logic;
			  input_zeros : in  STD_LOGIC_VECTOR (23 downto 0);
			  ENA_1 : IN  std_logic;
			  WEA_0 : IN  std_logic;
			  input1 : in  STD_LOGIC_VECTOR (7 downto 0);
			  input2 : in  STD_LOGIC_VECTOR (7 downto 0);
           output1 : out  STD_LOGIC_VECTOR (23 downto 0);
			  output2 : out  STD_LOGIC_VECTOR (23 downto 0)
			 );
end T_Box_2_port;

architecture T_Box_2_port_architecture of T_Box_2_port is

    type rom_type is array (0 to 255) of std_logic_vector (23 downto 0);                 
    signal ROM : rom_type:= ( X"C663A5",	
										X"F87C84",	
										X"EE7799",	
										X"F67B8D",	
										X"FFF20D",	
										X"D66BBD",	
										X"DE6FB1",	
										X"91C554",	
										X"603050",	
										X"020103",	
										X"CE67A9",	
										X"562B7D",	
										X"E7FE19",	
										X"B5D762",	
										X"4DABE6",	
										X"EC769A",	
										X"8FCA45",	
										X"1F829D",	
										X"89C940",	
										X"FA7D87",	
										X"EFFA15",	
										X"B259EB",	
										X"8E47C9",	
										X"FBF00B",	
										X"41ADEC",	
										X"B3D467",	
										X"5FA2FD",	
										X"45AFEA",	
										X"239CBF",	
										X"53A4F7",	
										X"E47296",	
										X"9BC05B",	
										X"75B7C2",	
										X"E1FD1C",	
										X"3D93AE",	
										X"4C266A",	
										X"6C365A",	
										X"7E3F41",	
										X"F5F702",	
										X"83CC4F",	
										X"68345C",	
										X"51A5F4",	
										X"D1E534",	
										X"F9F108",	
										X"E27193",	
										X"ABD873",	
										X"623153",	
										X"2A153F",	
										X"08040C",	
										X"95C752",	
										X"462365",	
										X"9DC35E",	
										X"301828",	
										X"3796A1",	
										X"0A050F",	
										X"2F9AB5",	
										X"0E0709",	
										X"241236",	
										X"1B809B",	
										X"DFE23D",	
										X"CDEB26",	
										X"4E2769",	
										X"7FB2CD",	
										X"EA759F",	
										X"12091B",	
										X"1D839E",	
										X"582C74",	
										X"341A2E",	
										X"361B2D",	
										X"DC6EB2",	
										X"B45AEE",	
										X"5BA0FB",	
										X"A452F6",	
										X"763B4D",	
										X"B7D661",	
										X"7DB3CE",	
										X"52297B",	
										X"DDE33E",	
										X"5E2F71",	
										X"138497",	
										X"A653F5",	
										X"B9D168",	
										X"000000",	
										X"C1ED2C",	
										X"402060",	
										X"E3FC1F",	
										X"79B1C8",	
										X"B65BED",	
										X"D46ABE",	
										X"8DCB46",	
										X"67BED9",	
										X"72394B",	
										X"944ADE",	
										X"984CD4",	
										X"B058E8",	
										X"85CF4A",	
										X"BBD06B",	
										X"C5EF2A",	
										X"4FAAE5",	
										X"EDFB16",	
										X"8643C5",	
										X"9A4DD7",	
										X"663355",	
										X"118594",	
										X"8A45CF",	
										X"E9F910",	
										X"040206",	
										X"FE7F81",	
										X"A050F0",	
										X"783C44",	
										X"259FBA",	
										X"4BA8E3",	
										X"A251F3",	
										X"5DA3FE",	
										X"8040C0",	
										X"058F8A",	
										X"3F92AD",	
										X"219DBC",	
										X"703848",	
										X"F1F504",	
										X"63BCDF",	
										X"77B6C1",	
										X"AFDA75",	
										X"422163",	
										X"201030",	
										X"E5FF1A",	
										X"FDF30E",	
										X"BFD26D",	
										X"81CD4C",	
										X"180C14",	
										X"261335",	
										X"C3EC2F",	
										X"BE5FE1",	
										X"3597A2",	
										X"8844CC",	
										X"2E1739",	
										X"93C457",	
										X"55A7F2",	
										X"FC7E82",	
										X"7A3D47",	
										X"C864AC",	
										X"BA5DE7",	
										X"32192B",	
										X"E67395",	
										X"C060A0",	
										X"198198",	
										X"9E4FD1",	
										X"A3DC7F",	
										X"442266",	
										X"542A7E",	
										X"3B90AB",	
										X"0B8883",	
										X"8C46CA",	
										X"C7EE29",	
										X"6BB8D3",	
										X"28143C",	
										X"A7DE79",	
										X"BC5EE2",	
										X"160B1D",	
										X"ADDB76",	
										X"DBE03B",	
										X"643256",	
										X"743A4E",	
										X"140A1E",	
										X"9249DB",	
										X"0C060A",	
										X"48246C",	
										X"B85CE4",	
										X"9FC25D",	
										X"BDD36E",	
										X"43ACEF",	
										X"C462A6",	
										X"3991A8",	
										X"3195A4",	
										X"D3E437",	
										X"F2798B",	
										X"D5E732",	
										X"8BC843",	
										X"6E3759",	
										X"DA6DB7",	
										X"018D8C",	
										X"B1D564",	
										X"9C4ED2",	
										X"49A9E0",	
										X"D86CB4",	
										X"AC56FA",	
										X"F3F407",	
										X"CFEA25",	
										X"CA65AF",	
										X"F47A8E",	
										X"47AEE9",	
										X"100818",	
										X"6FBAD5",	
										X"F07888",	
										X"4A256F",	
										X"5C2E72",	
										X"381C24",	
										X"57A6F1",	
										X"73B4C7",	
										X"97C651",	
										X"CBE823",	
										X"A1DD7C",	
										X"E8749C",	
										X"3E1F21",	
										X"964BDD",	
										X"61BDDC",	
										X"0D8B86",	
										X"0F8A85",	
										X"E07090",	
										X"7C3E42",	
										X"71B5C4",	
										X"CC66AA",	
										X"9048D8",	
										X"060305",	
										X"F7F601",	
										X"1C0E12",	
										X"C261A3",	
										X"6A355F",	
										X"AE57F9",	
										X"69B9D0",	
										X"178691",	
										X"99C158",	
										X"3A1D27",	
										X"279EB9",	
										X"D9E138",	
										X"EBF813",	
										X"2B98B3",	
										X"221133",	
										X"D269BB",	
										X"A9D970",	
										X"078E89",	
										X"3394A7",	
										X"2D9BB6",	
										X"3C1E22",	
										X"158792",	
										X"C9E920",	
										X"87CE49",	
										X"AA55FF",	
										X"502878",	
										X"A5DF7A",	
										X"038C8F",	
										X"59A1F8",	
										X"098980",	
										X"1A0D17",	
										X"65BFDA",	
										X"D7E631",	
										X"8442C6",	
										X"D068B8",	
										X"8241C3",	
										X"2999B0",	
										X"5A2D77",	
										X"1E0F11",	
										X"7BB0CB",	
										X"A854FC",	
										X"6DBBD6",	
										X"2C163A" );						  

begin

process (CLK)
begin
   if (CLK'event and CLK = '1') then
	
      if (ENA_1 = '1') then
		
         if (WEA_0 = '1') then
			
            ROM(conv_integer(input1)) <= input_zeros;
				
         end if;
			
			output1 <= ROM(conv_integer(input1));
			output2 <= ROM(conv_integer(input2));
		
      end if;
		
   end if;
	
end process;		

end T_Box_2_port_architecture;