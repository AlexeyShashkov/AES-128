library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity T_Box is
    port ( input : in  STD_LOGIC_VECTOR (7 downto 0);
           output : out  STD_LOGIC_VECTOR (23 downto 0)
			 );
end T_Box;

architecture T_Box_architecture of T_Box is

begin

	substitute: process(input)	
	begin
	
		case input is

			when X"00" => output <= X"C663A5";	
			when X"01" => output <= X"F87C84";	
			when X"02" => output <= X"EE7799";	
			when X"03" => output <= X"F67B8D";	
			when X"04" => output <= X"FFF20D";	
			when X"05" => output <= X"D66BBD";	
			when X"06" => output <= X"DE6FB1";	
			when X"07" => output <= X"91C554";	
			when X"08" => output <= X"603050";	
			when X"09" => output <= X"020103";	
			when X"0A" => output <= X"CE67A9";	
			when X"0B" => output <= X"562B7D";	
			when X"0C" => output <= X"E7FE19";	
			when X"0D" => output <= X"B5D762";	
			when X"0E" => output <= X"4DABE6";	
			when X"0F" => output <= X"EC769A";	
			when X"10" => output <= X"8FCA45";	
			when X"11" => output <= X"1F829D";	
			when X"12" => output <= X"89C940";	
			when X"13" => output <= X"FA7D87";	
			when X"14" => output <= X"EFFA15";	
			when X"15" => output <= X"B259EB";	
			when X"16" => output <= X"8E47C9";	
			when X"17" => output <= X"FBF00B";	
			when X"18" => output <= X"41ADEC";	
			when X"19" => output <= X"B3D467";	
			when X"1A" => output <= X"5FA2FD";	
			when X"1B" => output <= X"45AFEA";	
			when X"1C" => output <= X"239CBF";	
			when X"1D" => output <= X"53A4F7";	
			when X"1E" => output <= X"E47296";	
			when X"1F" => output <= X"9BC05B";	
			when X"20" => output <= X"75B7C2";	
			when X"21" => output <= X"E1FD1C";	
			when X"22" => output <= X"3D93AE";	
			when X"23" => output <= X"4C266A";	
			when X"24" => output <= X"6C365A";	
			when X"25" => output <= X"7E3F41";	
			when X"26" => output <= X"F5F702";	
			when X"27" => output <= X"83CC4F";	
			when X"28" => output <= X"68345C";	
			when X"29" => output <= X"51A5F4";	
			when X"2A" => output <= X"D1E534";	
			when X"2B" => output <= X"F9F108";	
			when X"2C" => output <= X"E27193";	
			when X"2D" => output <= X"ABD873";	
			when X"2E" => output <= X"623153";	
			when X"2F" => output <= X"2A153F";	
			when X"30" => output <= X"08040C";	
			when X"31" => output <= X"95C752";	
			when X"32" => output <= X"462365";	
			when X"33" => output <= X"9DC35E";	
			when X"34" => output <= X"301828";	
			when X"35" => output <= X"3796A1";	
			when X"36" => output <= X"0A050F";	
			when X"37" => output <= X"2F9AB5";	
			when X"38" => output <= X"0E0709";	
			when X"39" => output <= X"241236";	
			when X"3A" => output <= X"1B809B";	
			when X"3B" => output <= X"DFE23D";	
			when X"3C" => output <= X"CDEB26";	
			when X"3D" => output <= X"4E2769";	
			when X"3E" => output <= X"7FB2CD";	
			when X"3F" => output <= X"EA759F";	
			when X"40" => output <= X"12091B";	
			when X"41" => output <= X"1D839E";	
			when X"42" => output <= X"582C74";	
			when X"43" => output <= X"341A2E";	
			when X"44" => output <= X"361B2D";	
			when X"45" => output <= X"DC6EB2";	
			when X"46" => output <= X"B45AEE";	
			when X"47" => output <= X"5BA0FB";	
			when X"48" => output <= X"A452F6";	
			when X"49" => output <= X"763B4D";	
			when X"4A" => output <= X"B7D661";	
			when X"4B" => output <= X"7DB3CE";	
			when X"4C" => output <= X"52297B";	
			when X"4D" => output <= X"DDE33E";	
			when X"4E" => output <= X"5E2F71";	
			when X"4F" => output <= X"138497";	
			when X"50" => output <= X"A653F5";	
			when X"51" => output <= X"B9D168";	
			when X"52" => output <= X"000000";	
			when X"53" => output <= X"C1ED2C";	
			when X"54" => output <= X"402060";	
			when X"55" => output <= X"E3FC1F";	
			when X"56" => output <= X"79B1C8";	
			when X"57" => output <= X"B65BED";	
			when X"58" => output <= X"D46ABE";	
			when X"59" => output <= X"8DCB46";	
			when X"5A" => output <= X"67BED9";	
			when X"5B" => output <= X"72394B";	
			when X"5C" => output <= X"944ADE";	
			when X"5D" => output <= X"984CD4";	
			when X"5E" => output <= X"B058E8";	
			when X"5F" => output <= X"85CF4A";	
			when X"60" => output <= X"BBD06B";	
			when X"61" => output <= X"C5EF2A";	
			when X"62" => output <= X"4FAAE5";	
			when X"63" => output <= X"EDFB16";	
			when X"64" => output <= X"8643C5";	
			when X"65" => output <= X"9A4DD7";	
			when X"66" => output <= X"663355";	
			when X"67" => output <= X"118594";	
			when X"68" => output <= X"8A45CF";	
			when X"69" => output <= X"E9F910";	
			when X"6A" => output <= X"040206";	
			when X"6B" => output <= X"FE7F81";	
			when X"6C" => output <= X"A050F0";	
			when X"6D" => output <= X"783C44";	
			when X"6E" => output <= X"259FBA";	
			when X"6F" => output <= X"4BA8E3";	
			when X"70" => output <= X"A251F3";	
			when X"71" => output <= X"5DA3FE";	
			when X"72" => output <= X"8040C0";	
			when X"73" => output <= X"058F8A";	
			when X"74" => output <= X"3F92AD";	
			when X"75" => output <= X"219DBC";	
			when X"76" => output <= X"703848";	
			when X"77" => output <= X"F1F504";	
			when X"78" => output <= X"63BCDF";	
			when X"79" => output <= X"77B6C1";	
			when X"7A" => output <= X"AFDA75";	
			when X"7B" => output <= X"422163";	
			when X"7C" => output <= X"201030";	
			when X"7D" => output <= X"E5FF1A";	
			when X"7E" => output <= X"FDF30E";	
			when X"7F" => output <= X"BFD26D";	
			when X"80" => output <= X"81CD4C";	
			when X"81" => output <= X"180C14";	
			when X"82" => output <= X"261335";	
			when X"83" => output <= X"C3EC2F";	
			when X"84" => output <= X"BE5FE1";	
			when X"85" => output <= X"3597A2";	
			when X"86" => output <= X"8844CC";	
			when X"87" => output <= X"2E1739";	
			when X"88" => output <= X"93C457";	
			when X"89" => output <= X"55A7F2";	
			when X"8A" => output <= X"FC7E82";	
			when X"8B" => output <= X"7A3D47";	
			when X"8C" => output <= X"C864AC";	
			when X"8D" => output <= X"BA5DE7";	
			when X"8E" => output <= X"32192B";	
			when X"8F" => output <= X"E67395";	
			when X"90" => output <= X"C060A0";	
			when X"91" => output <= X"198198";	
			when X"92" => output <= X"9E4FD1";	
			when X"93" => output <= X"A3DC7F";	
			when X"94" => output <= X"442266";	
			when X"95" => output <= X"542A7E";	
			when X"96" => output <= X"3B90AB";	
			when X"97" => output <= X"0B8883";	
			when X"98" => output <= X"8C46CA";	
			when X"99" => output <= X"C7EE29";	
			when X"9A" => output <= X"6BB8D3";	
			when X"9B" => output <= X"28143C";	
			when X"9C" => output <= X"A7DE79";	
			when X"9D" => output <= X"BC5EE2";	
			when X"9E" => output <= X"160B1D";	
			when X"9F" => output <= X"ADDB76";	
			when X"A0" => output <= X"DBE03B";	
			when X"A1" => output <= X"643256";	
			when X"A2" => output <= X"743A4E";	
			when X"A3" => output <= X"140A1E";	
			when X"A4" => output <= X"9249DB";	
			when X"A5" => output <= X"0C060A";	
			when X"A6" => output <= X"48246C";	
			when X"A7" => output <= X"B85CE4";	
			when X"A8" => output <= X"9FC25D";	
			when X"A9" => output <= X"BDD36E";	
			when X"AA" => output <= X"43ACEF";	
			when X"AB" => output <= X"C462A6";	
			when X"AC" => output <= X"3991A8";	
			when X"AD" => output <= X"3195A4";	
			when X"AE" => output <= X"D3E437";	
			when X"AF" => output <= X"F2798B";	
			when X"B0" => output <= X"D5E732";	
			when X"B1" => output <= X"8BC843";	
			when X"B2" => output <= X"6E3759";	
			when X"B3" => output <= X"DA6DB7";	
			when X"B4" => output <= X"018D8C";	
			when X"B5" => output <= X"B1D564";	
			when X"B6" => output <= X"9C4ED2";	
			when X"B7" => output <= X"49A9E0";	
			when X"B8" => output <= X"D86CB4";	
			when X"B9" => output <= X"AC56FA";	
			when X"BA" => output <= X"F3F407";	
			when X"BB" => output <= X"CFEA25";	
			when X"BC" => output <= X"CA65AF";	
			when X"BD" => output <= X"F47A8E";	
			when X"BE" => output <= X"47AEE9";	
			when X"BF" => output <= X"100818";	
			when X"C0" => output <= X"6FBAD5";	
			when X"C1" => output <= X"F07888";	
			when X"C2" => output <= X"4A256F";	
			when X"C3" => output <= X"5C2E72";	
			when X"C4" => output <= X"381C24";	
			when X"C5" => output <= X"57A6F1";	
			when X"C6" => output <= X"73B4C7";	
			when X"C7" => output <= X"97C651";	
			when X"C8" => output <= X"CBE823";	
			when X"C9" => output <= X"A1DD7C";	
			when X"CA" => output <= X"E8749C";	
			when X"CB" => output <= X"3E1F21";	
			when X"CC" => output <= X"964BDD";	
			when X"CD" => output <= X"61BDDC";	
			when X"CE" => output <= X"0D8B86";	
			when X"CF" => output <= X"0F8A85";	
			when X"D0" => output <= X"E07090";	
			when X"D1" => output <= X"7C3E42";	
			when X"D2" => output <= X"71B5C4";	
			when X"D3" => output <= X"CC66AA";	
			when X"D4" => output <= X"9048D8";	
			when X"D5" => output <= X"060305";	
			when X"D6" => output <= X"F7F601";	
			when X"D7" => output <= X"1C0E12";	
			when X"D8" => output <= X"C261A3";	
			when X"D9" => output <= X"6A355F";	
			when X"DA" => output <= X"AE57F9";	
			when X"DB" => output <= X"69B9D0";	
			when X"DC" => output <= X"178691";	
			when X"DD" => output <= X"99C158";	
			when X"DE" => output <= X"3A1D27";	
			when X"DF" => output <= X"279EB9";	
			when X"E0" => output <= X"D9E138";	
			when X"E1" => output <= X"EBF813";	
			when X"E2" => output <= X"2B98B3";	
			when X"E3" => output <= X"221133";	
			when X"E4" => output <= X"D269BB";	
			when X"E5" => output <= X"A9D970";	
			when X"E6" => output <= X"078E89";	
			when X"E7" => output <= X"3394A7";	
			when X"E8" => output <= X"2D9BB6";	
			when X"E9" => output <= X"3C1E22";	
			when X"EA" => output <= X"158792";	
			when X"EB" => output <= X"C9E920";	
			when X"EC" => output <= X"87CE49";	
			when X"ED" => output <= X"AA55FF";	
			when X"EE" => output <= X"502878";	
			when X"EF" => output <= X"A5DF7A";	
			when X"F0" => output <= X"038C8F";	
			when X"F1" => output <= X"59A1F8";	
			when X"F2" => output <= X"098980";	
			when X"F3" => output <= X"1A0D17";	
			when X"F4" => output <= X"65BFDA";	
			when X"F5" => output <= X"D7E631";	
			when X"F6" => output <= X"8442C6";	
			when X"F7" => output <= X"D068B8";	
			when X"F8" => output <= X"8241C3";	
			when X"F9" => output <= X"2999B0";	
			when X"FA" => output <= X"5A2D77";	
			when X"FB" => output <= X"1E0F11";	
			when X"FC" => output <= X"7BB0CB";	
			when X"FD" => output <= X"A854FC";	
			when X"FE" => output <= X"6DBBD6";	
			when X"FF" => output <= X"2C163A";	 
			
			when others => null;
			
		end case;
		
	end process;

end T_Box_architecture;